`ifndef _GLB_MACROS_VH_
`define _GLB_MACROS_VH_

`define WORD_EXT(in_width, out_width, var) {{(out_width-in_width){1'b0}},var}

`endif