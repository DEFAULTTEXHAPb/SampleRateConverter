`ifndef _CTRL_VH_
`define _CTRL_VH_
`endif