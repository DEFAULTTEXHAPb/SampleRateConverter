`define VCC 1'b1
`define GND 1'b0