//! @title Coefficient address counter
//! @brief Counter for coefficient address
//! If `load` flag is active-high `coef_addr`
//! is set with value `coef_ptr` for coeffi-
//! cient downloading from CPU

module ctrl_ramdrv_coefcnt #(
    parameter integer ADDR_WIDTH = 12
) (
    input  wire                  clk,      //! __Clock__
    input  wire                  rst_n,      //! __Reset__
    input  wire                  load,     //! Coefficient load flag (and initial counter value set flag)
    input  wire                  cnt,      //! Counting enable
    input  wire [ADDR_WIDTH-1:0] coef_ptr, //! Initial coefficient pointer
    output wire [ADDR_WIDTH-1:0] coef_addr //! Output coefficient address
);
    
    //! Counter register
    reg [ADDR_WIDTH-1:0] coef_cnt = {ADDR_WIDTH{1'b0}};
    //! First cell address flag register
    reg                   first_register = 1'b1;

    assign coef_addr = coef_cnt;

    //! Counting process with counter value set
    always @(negedge clk) begin : coef_offset_counting
      if (rst_n == 1'b0) begin
        coef_cnt <= {ADDR_WIDTH{1'b0}};
        first_register <= 1'b1;
      end else if (load == 1'b1) begin
        coef_cnt <= coef_ptr;
        first_register <= 1'b1;
      end if (cnt == 1'b1) begin
        if (first_register == 1'b1) begin
          coef_cnt <= coef_cnt;
          first_register <= 1'b0;
        end else begin
          coef_cnt <= coef_cnt + 1'b1;          
        end
      end
    end

endmodule