`define DATA_PTR_W 12
`define MAX_STAGES     6
`define HEADER_PTR_WIDTH $clog2(64)